// uvm_sequencer的作用：
// 启动 sequence
// 将  sequence产生的item发送到UVM组件中(driver中)

// uvm_sequencer是拓展来的   #(my_transation)表示参数化的类
typedef uvm_sequencer #(my_transcation) my_sequencer; 


